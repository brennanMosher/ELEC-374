module NOT_FF(
 input [31:0] BusMuxOut,
 output Not_out);

endmodule 